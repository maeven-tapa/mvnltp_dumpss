module sample1 (A,B);
    input A;
    output B;
    assign B = A;

endmodule